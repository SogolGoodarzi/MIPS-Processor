module adder (a,b,s);
    input [31:0] a,b;
    output [31:0] s;
    assign s=a+b;
endmodule